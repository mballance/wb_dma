/****************************************************************************
 * dma_arb_agent_pkg.sv
 ****************************************************************************/

/**
 * Package: dma_arb_agent_pkg
 * 
 * TODO: Add package documentation
 */
package dma_arb_agent_pkg;
	`include "dma_arb_agent.svh"


endpackage


