/****************************************************************************
 * dma_config_pkg.sv
 ****************************************************************************/
 
`include "uvm_macros.svh"

/**
 * Package: dma_config_pkg
 * 
 * TODO: Add package documentation
 */
package dma_config_pkg;
	import uvm_pkg::*;
	import dma_reg_pkg::*;

	`include "dma_config_seq.svh"

endpackage


