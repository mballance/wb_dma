/****************************************************************************
 * memory_mgr_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: memory_mgr_pkg
 * 
 * TODO: Add package documentation
 */
package memory_mgr_pkg;
	import uvm_pkg::*;
	import wb_vip_pkg::*;

	`include "mem_ev.svh"
	`include "memory_mgr.svh"


endpackage


