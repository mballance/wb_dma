/****************************************************************************
 * dma_channel_reg.svh
 ****************************************************************************/

/**
 * Class: dma_channel_reg
 * 
 * TODO: Add class documentation
 */
class dma_channel_reg extends uvm_reg_block;
	`uvm_object_utils(dma_channel_reg)

	function new(string name="dma_channel_reg");

	endfunction


endclass


