/****************************************************************************
 * dma_arb_agent.svh
 ****************************************************************************/

/**
 * Class: dma_arb_agent
 * 
 * TODO: Add class documentation
 */
class dma_arb_agent extends uvm_agent;

	function new();

	endfunction


endclass


