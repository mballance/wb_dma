/****************************************************************************
 * dma_arb_config.svh
 ****************************************************************************/

/**
 * Class: dma_arb_config
 * 
 * TODO: Add class documentation
 */
class dma_arb_config extends uvm_sequence_item;

	function new();

	endfunction


endclass


