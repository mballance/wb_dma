/****************************************************************************
 * wb_dma_tests_pkg.sv
 ****************************************************************************/

/**
 * Package: wb_dma_tests_pkg
 * 
 * TODO: Add package documentation
 */
`include "uvm_macros.svh"
package wb_dma_tests_pkg;
	import uvm_pkg::*;
	import wb_dma_tb_pkg::*;
	
	`include "wb_dma_test_base.svh"


endpackage


