/****************************************************************************
 * dma_reg_pkg.sv
 ****************************************************************************/

/**
 * Package: dma_reg_pkg
 * 
 * TODO: Add package documentation
 */
package dma_reg_pkg;
	


endpackage


