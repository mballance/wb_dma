/****************************************************************************
 * timer_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: timer_pkg
 * 
 * TODO: Add package documentation
 */
package timer_pkg;
	import uvm_pkg::*;
	import wb_vip_pkg::*;

	`include "timer.svh"

endpackage


